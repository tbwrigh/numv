module numv

pub fn zero() int {
	return 0
}